module spi_dac (
    input clk100mhz,
    output reg cs,
    output reg mosi,
    output reg sclk,
    input st_wrt,
    input [11:0] data_in,
    output reg done
);

typedef enum logic [1:0] {idle_dac = 0, init_dac = 1, dac_data = 2, send_data = 3} state_type;
state_type state;

// Counter for DAC's output
integer count = 0;
reg [31:0] data = 32'h0;
reg [31:0] setup_dac = 32'h08000001;
reg dac_init = 1'b0;

// Local clock signals
integer clkdiv = 0;
reg clk1mhz = 1'b0;




// Clock generation process
always @(posedge clk100mhz) begin
    if (clkdiv == 49) 
    begin
        clkdiv <= 0;
        clk1mhz <= ~clk1mhz;
    end 
    else
    begin
        clkdiv <= clkdiv + 1;
    end
end

// DAC main process
always @(posedge clk1mhz or negedge st_wrt) begin
    if (!st_wrt) begin
        state <= idle_dac;
        cs    <= 1'b1;
        mosi  <= 1'b0;
        count <= 0;
        done <= 1'b0;
    end else begin
        case (state)
            idle_dac:
                begin
                    cs    <= 1'b1;
                    mosi  <= 1'b0;
                    count <= 0;
                    done  <= 1'b0;
                    if (!dac_init) 
                    begin
                        cs <= 1'b1;
                        state <= init_dac;
                    end 
                    else 
                    begin
                        cs <= 1'b1;
                        state <= dac_data;
                    end
                end
         
         //////////////////////initialize DAC to magic number
          
              init_dac : begin
               if(count < 32 )
                  begin
                  cs    <= 1'b0;
                  count <= count + 1;
                  mosi  <= setup_dac[31-count];
                  state <= init_dac;
                  end
               else
                 begin
                 count <= 0;
                 dac_init <= 1'b1;
                 cs <= 1'b1;
                 state <= dac_data;
                 end
              end
              
              		
					
              dac_data: begin
               cs   <= 1'b1;
               mosi <= 1'b0;
               data <= {12'h030, data_in, 8'h00 };
               state <= send_data;
              end
              
              send_data:
              begin
              if(count < 32)
                  begin
                  cs    <= 1'b0;
                  count <= count + 1;
                  mosi  <= data[31-count];
                  state <= send_data;
                  end
               else
                 begin
                 count    <= 0;
                 done     <= 1'b1;
                 cs       <= 1'b1;
                 state    <= idle_dac;
                 end
              end
          
          
            default:state <= idle_dac;
            
            
        endcase
    end
end

assign sclk = clk1mhz; // Drive DAC with locally generated 1MHz clock


endmodule

//////////////////////////////////////////////////////////

module tb_1;

    reg clk100mhz = 0;
    wire cs;
    wire mosi;
    wire sclk;
    reg st_wrt = 0;
    reg [11:0] data_in = 0;
    wire done;
    
    
    spi_dac dut (clk100mhz, cs, mosi, sclk, st_wrt, data_in, done);
    
    always#5 clk100mhz = ~clk100mhz;
    
    initial begin
    st_wrt = 1;
    data_in = 12'b101010101010;
    end



endmodule
